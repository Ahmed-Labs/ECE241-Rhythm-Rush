





module main()


//

parameter RED = 8'b2323423;
parameter BLUE = 8'b0234320;
parameter WHITE = 8'b0;





reg [10:0] score;
// score display

	reg [3:0] dig_2;
	reg [3:0] dig_1;
	reg [3:0] dig_0;


    

endmodule


module drawbox()
    input [2:0] colour_input;

endmodule