

module rythm_rush(

)

KEY 0-3: pressed 1-4
switch: 
    0 -> mouse click

endmodule